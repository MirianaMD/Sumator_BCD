module Sumator_tb#(parameter k=16);
  reg [k-1:0] x,y;
  wire [k:0] o;
  
  BCDp legat (.x(x), .y(y), .o(o));
	
	initial begin
	  
	 
	 /*
	 //8 biti
	 
	 
//37+89=126
#2 x=7'b00110111;
   y=7'b10001001;
#10 if(o==8'b100100110)
  $display("merge: %d %d %d",o[8],o[7:4],o[3:0]);
else   
  $display("nu merge: %d %d %d",o[8],o[7:4],o[3:0]);
  */
  
  
  
  
  //16 biti
  
  
//378+689=1067
#2 x=16'b0000001101111000;
   y=16'b0000011010001001;
#10 if(o==17'b00001000001100111)
  $display("merge: %d %d %d %d %d",o[16], o[15:12],o[11:8],o[7:4],o[3:0]);
else   
  $display("nu merge: %d %d %d %d %d",o[16], o[15:12],o[11:8],o[7:4],o[3:0]);
  
//437+578=1015
x=16'b0000010000110111;
y=16'b0000010101111000;
#10 if(o==17'b00001000000010101)
  $display("merge: %d %d %d %d %d",o[16], o[15:12],o[11:8],o[7:4],o[3:0]);
else   
  $display("nu merge: %d %d %d %d %d",o[16], o[15:12],o[11:8],o[7:4],o[3:0]);

//428+377=805
#2 x=15'b0000010000101000;
   y=15'b0000001101110111;
#10 if(o==16'b00000100000000101)
  $display("merge: %d %d %d %d %d",o[16], o[15:12],o[11:8],o[7:4],o[3:0]);
else   
  $display("nu merge: %d %d %d %d %d",o[16], o[15:12],o[11:8],o[7:4],o[3:0]);
  
//889+312=1201
#2 x=16'b0000100010001001;
   y=16'b0000001100010010;
#10 if(o==17'b00001001000000001)
  $display("merge: %d %d %d %d %d",o[16], o[15:12],o[11:8],o[7:4],o[3:0]);
else   
  $display("nu merge: %d %d %d %d %d",o[16], o[15:12],o[11:8],o[7:4],o[3:0]);

//888+312=1200//asta nu trebuia sa mearga intentionat
#2 x=16'b0000100010001000;
   y=16'b0000001100010010;
#10 if(o==17'b00001001000000001)
  $display("merge: %d %d %d %d %d",o[16], o[15:12],o[11:8],o[7:4],o[3:0]);
else   
  $display("nu merge: %d %d %d %d %d",o[16], o[15:12],o[11:8],o[7:4],o[3:0]);

//587+578=1165
x=16'b0000010110000111;
y=16'b0000010101111000;
#10 if(o==17'b00001000101100101)
  $display("merge: %d %d %d %d %d",o[16], o[15:12],o[11:8],o[7:4],o[3:0]);
else   
  $display("nu merge: %d %d %d %d %d",o[16], o[15:12],o[11:8],o[7:4],o[3:0]);

//1587+578=2165
x=16'b0001010110000111;
y=16'b0000010101111000;
#10 if(o==17'b00010000101100101)
  $display("merge: %d %d %d %d %d",o[16], o[15:12],o[11:8],o[7:4],o[3:0]);
else   
  $display("nu merge: %d %d %d %d %d",o[16], o[15:12],o[11:8],o[7:4],o[3:0]);

//33+33=66
x=16'b0000000000110011;
y=16'b0000000000110011;
#10 if(o==17'b00000000001100110)
  $display("merge: %d %d %d %d %d",o[16], o[15:12],o[11:8],o[7:4],o[3:0]);
else   
  $display("nu merge: %d %d %d %d %d",o[16], o[15:12],o[11:8],o[7:4],o[3:0]);

//0+66=66
x=16'b0000000000000000;
y=16'b0000000001100110;
#10 if(o==17'b00000000001100110)
  $display("merge: %d %d %d %d %d",o[16], o[15:12],o[11:8],o[7:4],o[3:0]);
else   
  $display("nu merge: %d %d %d %d %d",o[16], o[15:12],o[11:8],o[7:4],o[3:0]);
  
//9999+7779=17778
x=16'b1001100110011001;
y=16'b0111011101111001;
#10 if(o==17'b10111011101111000)
  $display("merge: %d %d %d %d %d",o[16], o[15:12],o[11:8],o[7:4],o[3:0]);
else   
  $display("nu merge: %d %d %d %d %d",o[16], o[15:12],o[11:8],o[7:4],o[3:0]);
  
  
  
  /*
  //32 de biti
  
  
  
//17778+99999=117777;
x=31'b00000000000000010111011101111000;
y=31'b00000000000010011001100110011001;
#10 if(o==32'b00000000000100010111011101110111)
  $display("merge: %d %d %d %d %d %d %d %d %d",o[32], o[31:28], o[27:24], o[23:20], o[19:16], o[15:12], o[11:8], o[7:4], o[3:0]);
else   
  $display("nu merge: %d %d %d %d %d %d %d %d %d",o[32], o[31:28], o[27:24], o[23:20], o[19:16], o[15:12], o[11:8], o[7:4], o[3:0]);
*/

end
	
endmodule